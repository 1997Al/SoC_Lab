module zeroTruncBits(o_Out);
    output  o_Out;

    assign o_Out = 0;

endmodule
